--
--    Digits Box: takes in 3 digits (from 0 to 9) and prints those digits on the 
--                vga monitor.
--    
--    Module of:
--        - vga_module
--
--    Internal singals:
--        - sig_0 - sig_10: A 5x5 matrix that contains a digit from 0-9
--        - sig_dec: A matrix the contains an image of a decimal point
--        - box_loc_x/y_min/max: Min and max indices from x and y
--        - pixel_color: Colour of an individual pixel


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity digits_box is
    Port (
            clk:          in  STD_LOGIC;
            reset:        in  STD_LOGIC;

            distance_bcd: in  STD_LOGIC_VECTOR(4*4-1 downto 0);

            scan_line_x:  in  STD_LOGIC_VECTOR(10 downto 0);
            scan_line_y:  in  STD_LOGIC_VECTOR(10 downto 0);
            --kHz:          in  STD_LOGIC;
            red:          out STD_LOGIC_VECTOR(3 downto 0);
            blue:         out STD_LOGIC_VECTOR(3 downto 0);
            green:        out std_logic_vector(3 downto 0)
          );
end digits_box;

architecture Behavioral of digits_box is

-- Internal Signals  -----------------------------------------------------------
    type MAT is array (24 downto 0) of std_logic_vector(24 downto 0);
    constant sig_E: Mat := (("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"));
    constant sig_D: Mat := (("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"));
    constant sig_0: MAT := (("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"));
    constant sig_1: MAT := (("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"), ("0000000000000000000000000"));
    constant sig_2: MAT := (("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111111111000000000011111"), ("1111111111000000000011111"), ("1111111111000000000011111"), ("1111111111000000000011111"), ("1111111111000000000011111"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"));
    constant sig_3: MAT := (("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"));
    constant sig_4: MAT := (("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"));
    constant sig_5: MAT := (("1111111111000000000011111"), ("1111111111000000000011111"), ("1111111111000000000011111"), ("1111111111000000000011111"), ("1111111111000000000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000001111111111"), ("1111100000000001111111111"), ("1111100000000001111111111"), ("1111100000000001111111111"), ("1111100000000001111111111"));
    constant sig_6: MAT := (("0000011111000000000011111"), ("0000011111000000000011111"), ("0000011111000000000011111"), ("0000011111000000000011111"), ("0000011111000000000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"));
    constant sig_7: MAT := (("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000001111111111"), ("0000000000000001111111111"), ("0000000000000001111111111"), ("0000000000000001111111111"), ("0000000000000001111111111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000000000111110000011111"), ("0000011111000000000011111"), ("0000011111000000000011111"), ("0000011111000000000011111"), ("0000011111000000000011111"), ("0000011111000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"));
    constant sig_8: MAT := (("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"));
    constant sig_9: MAT := (("0000000000111111111111111"), ("0000000000111111111111111"), ("0000000000111111111111111"), ("0000000000111111111111111"), ("0000000000111111111111111"), ("0000011111111110000011111"), ("0000011111111110000011111"), ("0000011111111110000011111"), ("0000011111111110000011111"), ("0000011111111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000111110000011111"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"), ("1111100000000001111100000"));

    constant box_loc_x_min: STD_LOGIC_VECTOR(9 downto 0) := "0000000000";
    constant box_loc_y_min: STD_LOGIC_VECTOR(9 downto 0) := "0000000000";
    constant box_loc_x_max: STD_LOGIC_VECTOR(9 downto 0) := "1001111111"; -- 640-1 -- 640 is 1010000000
    constant box_loc_y_max: STD_LOGIC_VECTOR(9 downto 0) := "0111011111"; -- 480-1 -- 480 is 0111100000
    signal pixel_color:     STD_LOGIC_VECTOR(11 downto 0);
   
    signal current_digit_value: STD_LOGIC_VECTOR(3 downto 0); -- Value of the digit you are currently in (or 0s)
    signal output_digit: MAT;

    constant pos_start_x_sig_digit_d1:  STD_LOGIC_VECTOR(9 downto 0) := "0000010000"; -- 16
    constant pos_start_x_sig_digit_d2:  STD_LOGIC_VECTOR(9 downto 0) := "0000101101"; -- 45
    constant pos_start_x_sig_digit_d3:  STD_LOGIC_VECTOR(9 downto 0) := "0001001010"; -- 74
    constant pos_start_x_sig_digit_d4:  STD_LOGIC_VECTOR(9 downto 0) := "0001100111"; -- 103
    constant pos_end_x_sig_digit_d1:    STD_LOGIC_VECTOR(9 downto 0) := "0000101001"; -- 41
    constant pos_end_x_sig_digit_d2:    STD_LOGIC_VECTOR(9 downto 0) := "0001000110"; -- 70
    constant pos_end_x_sig_digit_d3:    STD_LOGIC_VECTOR(9 downto 0) := "0001100011"; -- 99
    constant pos_end_x_sig_digit_d4:    STD_LOGIC_VECTOR(9 downto 0) := "0010000000"; -- 128
    constant pos_start_y:               STD_LOGIC_VECTOR(9 downto 0) := "0000010000"; -- 16 -- All digits share these
    constant pos_end_y:                 STD_LOGIC_VECTOR(9 downto 0) := "0000101001"; -- 41 -- All digits share these

    signal currently_sig_digit_d1:      STD_LOGIC := '0';
    signal currently_sig_digit_d2:      STD_LOGIC := '0';
    signal currently_sig_digit_d4:      STD_LOGIC := '0';
    signal currently_sig_digit_d3:      STD_LOGIC := '0';
    signal pos_start_x_current_sig:     STD_LOGIC_VECTOR(9 downto 0); -- The pos_start_x_sig for the current digit
    signal current_sig_x_offset:        integer := 0; -- Used for indexing the current sig_digit MAT
    signal current_sig_y_offset:        integer := 0;

begin


-- Internal processes  ---------------------------------------------------------
    -- Figure out which digit (if any is currently being shown)
        currently_sig_digit_d1 <= '1'
                when (scan_line_x >= pos_start_x_sig_digit_d1) AND
                     (scan_line_x <  pos_end_x_sig_digit_d1) AND
                     (scan_line_y >= pos_start_y) AND
                     (scan_line_y <  pos_end_y) 
                else '0';
        currently_sig_digit_d2 <= '1'
                when (scan_line_x >= pos_start_x_sig_digit_d2) AND
                     (scan_line_x <  pos_end_x_sig_digit_d2) AND
                     (scan_line_y >= pos_start_y) AND
                     (scan_line_y <  pos_end_y) 
                else '0';
        currently_sig_digit_d3 <= '1'
                when (scan_line_x >= pos_start_x_sig_digit_d3) AND
                     (scan_line_x <  pos_end_x_sig_digit_d3) AND
                     (scan_line_y >= pos_start_y) AND
                     (scan_line_y <  pos_end_y) 
                else '0';
        currently_sig_digit_d4 <= '1'
                when (scan_line_x >= pos_start_x_sig_digit_d4) AND
                     (scan_line_x <  pos_end_x_sig_digit_d4) AND
                     (scan_line_y >= pos_start_y) AND
                     (scan_line_y <  pos_end_y) 
                else '0';

    -- Get the x & y offset INSIDE a digit
        -- The starting pos of the digit you are currently in (or 0s if not in digit)
        pos_start_x_current_sig <=   pos_start_x_sig_digit_d1 when (currently_sig_digit_d1 = '1')
                                else pos_start_x_sig_digit_d2 when (currently_sig_digit_d2 = '1')
                                else pos_start_x_sig_digit_d3 when (currently_sig_digit_d3 = '1')
                                else pos_start_x_sig_digit_d4 when (currently_sig_digit_d4 = '1')
                                else (others => '0');
        -- Determine how many pixels from the start of the current digit the scan lines are
        current_sig_x_offset <= CONV_INTEGER(UNSIGNED(scan_line_x - pos_start_x_current_sig));
        current_sig_y_offset <= CONV_INTEGER(UNSIGNED(scan_line_y - pos_start_y));

    -- Get the values of the current digits
        current_digit_value <=
                distance_bcd(4*4-1 downto 3*4) when (currently_sig_digit_d1 = '1')
                else distance_bcd(4*3-1 downto 2*4) when (currently_sig_digit_d2 = '1')
                else distance_bcd(4*2-1 downto 1*4) when (currently_sig_digit_d3 = '1')
                else distance_bcd(4*1-1 downto 0*4) when (currently_sig_digit_d4 = '1')
                else (others => '0');
 
        CURRENT_DIGIT: process(current_digit_value)
        begin
            case current_digit_value is
                when "0000" => output_digit <= sig_0;
                when "0001" => output_digit <= sig_1;
                when "0010" => output_digit <= sig_2;
                when "0011" => output_digit <= sig_3;
                when "0100" => output_digit <= sig_4;
                when "0101" => output_digit <= sig_5;
                when "0110" => output_digit <= sig_6;
                when "0111" => output_digit <= sig_7;
                when "1000" => output_digit <= sig_8;
                when "1001" => output_digit <= sig_9;
                when "1110" => output_digit <= sig_D;
                when others => output_digit <= sig_E;
            end case;
        end process;

    -- Select the color
        pixel_color <= "111011111111"
                  when  ((output_digit(current_sig_x_offset)(current_sig_y_offset) = '1')) AND 
                         ((currently_sig_digit_d1 = '1') OR
                         (currently_sig_digit_d2 = '1') OR
                         (currently_sig_digit_d4 = '1') OR
                         (currently_sig_digit_d3 = '1'))
                else
                         "000000000000"; -- represents background color

                                
red   <= pixel_color(11 downto 8);
green <= pixel_color(7 downto 4);
blue  <= pixel_color(3 downto 0);


end Behavioral;
