library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    use IEEE.STD_LOGIC_ARITH.ALL;
    use IEEE.STD_LOGIC_UNSIGNED.ALL;
    
    entity estimator is
            generic (width: integer := 9);
            Port (
                    clk        : in  STD_LOGIC;
                    reset      : in  STD_LOGIC;
                    en_dists_cm: in  STD_LOGIC;
                    en_dists_in: in  STD_LOGIC;
                    voltage    : in  STD_LOGIC_VECTOR(width-1 downto 0);
                    distance   : out STD_LOGIC_VECTOR(4*4-1 downto 0)
            );
    end estimator;
    
    architecture Behavioral of estimator is
    type ROM is array (0 to 511) of STD_LOGIC_VECTOR(4*4-1 downto 0);
    constant dists_cm: ROM := (("0111011111000110"), ("0111011011001000"), ("0111010111001001"), ("0111010111000001"), ("0111010011000011"), ("0111001111000101"), ("0111001011000111"), ("0111000111001001"), ("0111000111000001"), ("0111000011000011"), ("0110100111000101"), ("0110100011000111"), ("0110100011000000"), ("0110011111000010"), ("0110011011000101"), ("0110010111000111"), ("0110010111000000"), ("0110010011000011"), ("0110001111000101"), ("0110001011001000"), ("0110001011000001"), ("0110000111000100"), ("0110000011000111"), ("0110000011000001"), ("0101100111000100"), ("0101100011000111"), ("0101100011000001"), ("0101011111000100"), ("0101011011001000"), ("0101011011000001"), ("0101010111000101"), ("0101010011001000"), ("0101010011000010"), ("0101001111000110"), ("0101001111000000"), ("0101001011000100"), ("0101000111001000"), ("0101000111000010"), ("0101000011000110"), ("0101000011000000"), ("0100100111000101"), ("0100100011001001"), ("0100100011000011"), ("0100011111001000"), ("0100011111000010"), ("0100011011000111"), ("0100011011000010"), ("0100010111000110"), ("0100010111000001"), ("0100010011000110"), ("0100010011000001"), ("0100001111000110"), ("0100001111000001"), ("0100001011000110"), ("0100001011000001"), ("0100000111000110"), ("0100000111000001"), ("0100000011000110"), ("0100000011000010"), ("0011100111000111"), ("0011100111000011"), ("0011100011001000"), ("0011100011000100"), ("0011011111001001"), ("0011011111000101"), ("0011011111000000"), ("0011011011000110"), ("0011011011000010"), ("0011010111001000"), ("0011010111000100"), ("0011010111000000"), ("0011010011000110"), ("0011010011000010"), ("0011001111001000"), ("0011001111000100"), ("0011001111000000"), ("0011001011000110"), ("0011001011000010"), ("0011000111001001"), ("0011000111000101"), ("0011000111000001"), ("0011000011001000"), ("0011000011000100"), ("0011000011000001"), ("0010100111000111"), ("0010100111000100"), ("0010100111000001"), ("0010100011000111"), ("0010100011000100"), ("0010100011000001"), ("0010011111001000"), ("0010011111000100"), ("0010011111000001"), ("0010011011001000"), ("0010011011000101"), ("0010011011000010"), ("0010010111001001"), ("0010010111000110"), ("0010010111000011"), ("0010010111000001"), ("0010010011001000"), ("0010010011000101"), ("0010010011000010"), ("0010001111001001"), ("0010001111000111"), ("0010001111000100"), ("0010001111000010"), ("0010001011001001"), ("0010001011000111"), ("0010001011000100"), ("0010001011000010"), ("0010000111001001"), ("0010000111000111"), ("0010000111000100"), ("0010000111000010"), ("0010000111000000"), ("0010000011000111"), ("0010000011000101"), ("0010000011000011"), ("0010000011000001"), ("0001100111001001"), ("0001100111000111"), ("0001100111000101"), ("0001100111000010"), ("0001100111000000"), ("0001100011001000"), ("0001100011000110"), ("0001100011000101"), ("0001100011000011"), ("0001100011000001"), ("0001011111001001"), ("0001011111000111"), ("0001011111000101"), ("0001011111000011"), ("0001011111000010"), ("0001011111000000"), ("0001011011001000"), ("0001011011000111"), ("0001011011000101"), ("0001011011000011"), ("0001011011000010"), ("0001011011000000"), ("0001010111001001"), ("0001010111000111"), ("0001010111000101"), ("0001010111000100"), ("0001010111000011"), ("0001010111000001"), ("0001010111000000"), ("0001010011001000"), ("0001010011000111"), ("0001010011000101"), ("0001010011000100"), ("0001010011000011"), ("0001010011000010"), ("0001010011000000"), ("0001001111001001"), ("0001001111001000"), ("0001001111000111"), ("0001001111000101"), ("0001001111000100"), ("0001001111000011"), ("0001001111000010"), ("0001001111000001"), ("0001001111000000"), ("0001001011001000"), ("0001001011000111"), ("0001001011000110"), ("0001001011000101"), ("0001001011000100"), ("0001001011000011"), ("0001001011000010"), ("0001001011000001"), ("0001001011000000"), ("0001000111001001"), ("0001000111001000"), ("0001000111000111"), ("0001000111000111"), ("0001000111000110"), ("0001000111000101"), ("0001000111000100"), ("0001000111000011"), ("0001000111000010"), ("0001000111000001"), ("0001000111000001"), ("0001000111000000"), ("0001000011001001"), ("0001000011001000"), ("0001000011000111"), ("0001000011000111"), ("0001000011000110"), ("0001000011000101"), ("0001000011000100"), ("0001000011000100"), ("0001000011000011"), ("0001000011000010"), ("0001000011000010"), ("0001000011000001"), ("0001000011000000"), ("0001000011000000"), ("1001110010010110"), ("1001110010001001"), ("1001110010000011"), ("1001110001110111"), ("1001110001110001"), ("1001110001100101"), ("1001110001011001"), ("1001110001010100"), ("1001110001001000"), ("1001110001000010"), ("1001110000110111"), ("1001110000110001"), ("1001110000100110"), ("1001110000100001"), ("1001110000010110"), ("1001110000010001"), ("1001110000000110"), ("1001110000000001"), ("1000110010010110"), ("1000110010010001"), ("1000110010000110"), ("1000110010000001"), ("1000110001110111"), ("1000110001110010"), ("1000110001101000"), ("1000110001100011"), ("1000110001011001"), ("1000110001010100"), ("1000110001010000"), ("1000110001000110"), ("1000110001000001"), ("1000110000110111"), ("1000110000110011"), ("1000110000101001"), ("1000110000100101"), ("1000110000100001"), ("1000110000010111"), ("1000110000010011"), ("1000110000001001"), ("1000110000000101"), ("1000110000000001"), ("0111110010011000"), ("0111110010010100"), ("0111110010010000"), ("0111110010000111"), ("0111110010000011"), ("0111110001111001"), ("0111110001110110"), ("0111110001110010"), ("0111110001101001"), ("0111110001100101"), ("0111110001100010"), ("0111110001011000"), ("0111110001010101"), ("0111110001010001"), ("0111110001001000"), ("0111110001000101"), ("0111110001000001"), ("0111110000111000"), ("0111110000110101"), ("0111110000110001"), ("0111110000101000"), ("0111110000100101"), ("0111110000100001"), ("0111110000011000"), ("0111110000010101"), ("0111110000010010"), ("0111110000001001"), ("0111110000000101"), ("0111110000000010"), ("0110110010011001"), ("0110110010010110"), ("0110110010010011"), ("0110110010010000"), ("0110110010000110"), ("0110110010000011"), ("0110110010000000"), ("0110110001110111"), ("0110110001110100"), ("0110110001110001"), ("0110110001101000"), ("0110110001100101"), ("0110110001100001"), ("0110110001011000"), ("0110110001010101"), ("0110110001010010"), ("0110110001001001"), ("0110110001000110"), ("0110110001000011"), ("0110110001000000"), ("0110110000110111"), ("0110110000110011"), ("0110110000110000"), ("0110110000100111"), ("0110110000100100"), ("0110110000100001"), ("0110110000011000"), ("0110110000010101"), ("0110110000010010"), ("0110110000001000"), ("0110110000000101"), ("0110110000000010"), ("0101110010011001"), ("0101110010010110"), ("0101110010010011"), ("0101110010010000"), ("0101110010000111"), ("0101110010000011"), ("0101110010000000"), ("0101110001110111"), ("0101110001110100"), ("0101110001110001"), ("0101110001101000"), ("0101110001100100"), ("0101110001100001"), ("0101110001011000"), ("0101110001010101"), ("0101110001010010"), ("0101110001001001"), ("0101110001000101"), ("0101110001000010"), ("0101110000111001"), ("0101110000110110"), ("0101110000110011"), ("0101110000101001"), ("0101110000100110"), ("0101110000100011"), ("0101110000100000"), ("0101110000010111"), ("0101110000010011"), ("0101110000010000"), ("0101110000000111"), ("0101110000000100"), ("0101110000000001"), ("0100110010010111"), ("0100110010010100"), ("0100110010010001"), ("0100110010001000"), ("0100110010000101"), ("0100110010000010"), ("0100110001111000"), ("0100110001110101"), ("0100110001110010"), ("0100110001101001"), ("0100110001100110"), ("0100110001100011"), ("0100110001100000"), ("0100110001010111"), ("0100110001010011"), ("0100110001010000"), ("0100110001000111"), ("0100110001000100"), ("0100110001000001"), ("0100110000111000"), ("0100110000110101"), ("0100110000110010"), ("0100110000101001"), ("0100110000100110"), ("0100110000100011"), ("0100110000100000"), ("0100110000010111"), ("0100110000010100"), ("0100110000010010"), ("0100110000001001"), ("0100110000000110"), ("0100110000000011"), ("0100110000000000"), ("0011110010011000"), ("0011110010010101"), ("0011110010010010"), ("0011110010010000"), ("0011110010000111"), ("0011110010000100"), ("0011110010000010"), ("0011110001111001"), ("0011110001110111"), ("0011110001110100"), ("0011110001110010"), ("0011110001110000"), ("0011110001100111"), ("0011110001100101"), ("0011110001100011"), ("0011110001100000"), ("0011110001011000"), ("0011110001010110"), ("0011110001010100"), ("0011110001010010"), ("0011110001010000"), ("0011110001001000"), ("0011110001000110"), ("0011110001000100"), ("0011110001000011"), ("0011110001000001"), ("0011110000111001"), ("0011110000111000"), ("0011110000110110"), ("0011110000110101"), ("0011110000110011"), ("0011110000110010"), ("0011110000110001"), ("0011110000110000"), ("0011110000101001"), ("0011110000101000"), ("0011110000100111"), ("0011110000100110"), ("0011110000100101"), ("0011110000100100"), ("0011110000100011"), ("0011110000100011"), ("0011110000100010"), ("0011110000100010"), ("0011110000100010"), ("0011110000100001"), ("0011110000100001"), ("0011110000100001"), ("0011110000100001"), ("0011110000100010"), ("0011110000100010"), ("0011110000100010"), ("0011110000100011"), ("0011110000100011"), ("0011110000100100"), ("0011110000100101"), ("0011110000100101"), ("0011110000100110"), ("0011110000101000"), ("0011110000101001"), ("0011110000110000"), ("0011110000110010"), ("0011110000110011"), ("0011110000110101"), ("0011110000110111"), ("0011110000111001"), ("0011110001000001"), ("0011110001000011"), ("0011110001000110"), ("0011110001001000"), ("0011110001010001"), ("0011110001010011"), ("0011110001010110"), ("0011110001011001"), ("0011110001100011"), ("0011110001100110"), ("0011110001110000"), ("0011110001110011"), ("0011110001110111"), ("0011110010000001"), ("0011110010000101"), ("0011110010010000"), ("0011110010010100"), ("0011110010011001"), ("0100110000000100"), ("0100110000001001"), ("0100110000010100"), ("0100110000011001"), ("0100110000100101"), ("0100110000110001"), ("0100110000110111"), ("0100110001000011"), ("0100110001001001"), ("0100110001010110"), ("0100110001100010"), ("0100110001101001"), ("0100110001110110"), ("0100110010000100"), ("0100110010010001"), ("0100110010011001"), ("0101110000000111"), ("0101110000010101"), ("0101110000100100"), ("0101110000110010"), ("0101110001000001"), ("0101110001010000"), ("0101110001011001"), ("0101110001101001"), ("0101110001111001"), ("0101110010001001"), ("0101110010011001"), ("0110110000010000"), ("0110110000100000"), ("0110110000110001"), ("0110110001000011"), ("0110110001010100"), ("0110110001100110"), ("0110110001111000"), ("0110110010010000"), ("0111110000000011"), ("0111110000010110"), ("0111110000101001"), ("0111110001000010"), ("0111110001010110"), ("0111110001110000"), ("0111110010000100"), ("0111110010011001"), ("1000110000010100"), ("1000110000101001"), ("1000110001000100"), ("1000110001100000"), ("1000110001110110"), ("1000110010010010"), ("1001110000001001"), ("1001110000100110"), ("1001110001000011"), ("1001110001100001"), ("1001110001111001"), ("1001110010010111"), ("0001000011000001"), ("0001000011000011"), ("0001000011000101"), ("0001000011000111"), ("0001000011001001"), ("0001000111000001"));
    constant dists_in: ROM := (("0011000011000101"), ("0011000011000010"), ("0010100111001001"), ("0010100111000101"), ("0010100111000010"), ("0010100011001001"), ("0010100011000110"), ("0010100011000011"), ("0010011111001001"), ("0010011111000110"), ("0010011111000011"), ("0010011111000000"), ("0010011011000111"), ("0010011011000100"), ("0010011011000001"), ("0010010111001000"), ("0010010111000110"), ("0010010111000011"), ("0010010111000000"), ("0010010011000111"), ("0010010011000100"), ("0010010011000010"), ("0010001111001001"), ("0010001111000110"), ("0010001111000100"), ("0010001111000001"), ("0010001011001000"), ("0010001011000110"), ("0010001011000011"), ("0010001011000001"), ("0010000111001000"), ("0010000111000110"), ("0010000111000011"), ("0010000111000001"), ("0010000011001000"), ("0010000011000110"), ("0010000011000100"), ("0010000011000001"), ("0001100111001001"), ("0001100111000111"), ("0001100111000100"), ("0001100111000010"), ("0001100111000000"), ("0001100011001000"), ("0001100011000110"), ("0001100011000100"), ("0001100011000001"), ("0001011111001001"), ("0001011111000111"), ("0001011111000101"), ("0001011111000011"), ("0001011111000001"), ("0001011011001001"), ("0001011011000111"), ("0001011011000101"), ("0001011011000011"), ("0001011011000010"), ("0001011011000000"), ("0001010111001000"), ("0001010111000110"), ("0001010111000100"), ("0001010111000010"), ("0001010111000001"), ("0001010011001001"), ("0001010011000111"), ("0001010011000110"), ("0001010011000100"), ("0001010011000010"), ("0001010011000001"), ("0001001111001001"), ("0001001111000111"), ("0001001111000110"), ("0001001111000100"), ("0001001111000011"), ("0001001111000001"), ("0001001111000000"), ("0001001011001000"), ("0001001011000111"), ("0001001011000101"), ("0001001011000100"), ("0001001011000010"), ("0001001011000001"), ("0001000111001001"), ("0001000111001000"), ("0001000111000111"), ("0001000111000101"), ("0001000111000100"), ("0001000111000011"), ("0001000111000001"), ("0001000111000000"), ("0001000011001001"), ("0001000011001000"), ("0001000011000110"), ("0001000011000101"), ("0001000011000100"), ("0001000011000011"), ("0001000011000010"), ("0001000011000001"), ("1001110010011001"), ("1001110010001000"), ("1001110001110111"), ("1001110001100110"), ("1001110001010101"), ("1001110001000100"), ("1001110000110100"), ("1001110000100011"), ("1001110000010011"), ("1001110000000011"), ("1000110010010011"), ("1000110010000011"), ("1000110001110100"), ("1000110001100100"), ("1000110001010101"), ("1000110001000101"), ("1000110000110110"), ("1000110000100111"), ("1000110000011000"), ("1000110000010000"), ("1000110000000001"), ("0111110010010010"), ("0111110010000100"), ("0111110001110110"), ("0111110001100111"), ("0111110001011001"), ("0111110001010001"), ("0111110001000011"), ("0111110000110110"), ("0111110000101000"), ("0111110000100000"), ("0111110000010011"), ("0111110000000110"), ("0110110010011000"), ("0110110010010001"), ("0110110010000100"), ("0110110001110111"), ("0110110001110001"), ("0110110001100100"), ("0110110001010111"), ("0110110001010001"), ("0110110001000100"), ("0110110000111000"), ("0110110000110010"), ("0110110000100110"), ("0110110000100000"), ("0110110000010100"), ("0110110000001000"), ("0110110000000010"), ("0101110010010110"), ("0101110010010001"), ("0101110010000101"), ("0101110010000000"), ("0101110001110100"), ("0101110001101001"), ("0101110001100100"), ("0101110001011001"), ("0101110001010100"), ("0101110001001001"), ("0101110001000100"), ("0101110000111001"), ("0101110000110100"), ("0101110000101001"), ("0101110000100101"), ("0101110000100000"), ("0101110000010110"), ("0101110000010001"), ("0101110000000111"), ("0101110000000011"), ("0100110010011001"), ("0100110010010101"), ("0100110010010001"), ("0100110010000111"), ("0100110010000011"), ("0100110001111001"), ("0100110001110101"), ("0100110001110001"), ("0100110001100111"), ("0100110001100100"), ("0100110001100000"), ("0100110001010111"), ("0100110001010011"), ("0100110001010000"), ("0100110001000110"), ("0100110001000011"), ("0100110001000000"), ("0100110000110111"), ("0100110000110100"), ("0100110000110000"), ("0100110000100111"), ("0100110000100100"), ("0100110000100001"), ("0100110000011000"), ("0100110000010110"), ("0100110000010011"), ("0100110000010000"), ("0100110000000111"), ("0100110000000101"), ("0100110000000010"), ("0011110010011001"), ("0011110010010111"), ("0011110010010100"), ("0011110010010010"), ("0011110010001001"), ("0011110010000111"), ("0011110010000100"), ("0011110010000010"), ("0011110010000000"), ("0011110001110111"), ("0011110001110101"), ("0011110001110011"), ("0011110001110001"), ("0011110001101001"), ("0011110001100110"), ("0011110001100100"), ("0011110001100010"), ("0011110001100000"), ("0011110001011000"), ("0011110001010110"), ("0011110001010100"), ("0011110001010010"), ("0011110001010000"), ("0011110001001001"), ("0011110001000111"), ("0011110001000101"), ("0011110001000011"), ("0011110001000001"), ("0011110000111001"), ("0011110000111000"), ("0011110000110110"), ("0011110000110100"), ("0011110000110011"), ("0011110000110001"), ("0011110000101001"), ("0011110000101000"), ("0011110000100110"), ("0011110000100100"), ("0011110000100011"), ("0011110000100001"), ("0011110000100000"), ("0011110000011000"), ("0011110000010111"), ("0011110000010101"), ("0011110000010100"), ("0011110000010010"), ("0011110000010001"), ("0011110000001001"), ("0011110000001000"), ("0011110000000111"), ("0011110000000101"), ("0011110000000100"), ("0011110000000010"), ("0011110000000001"), ("0011110000000000"), ("0010110010011000"), ("0010110010010111"), ("0010110010010110"), ("0010110010010100"), ("0010110010010011"), ("0010110010010010"), ("0010110010010000"), ("0010110010001001"), ("0010110010001000"), ("0010110010000110"), ("0010110010000101"), ("0010110010000100"), ("0010110010000010"), ("0010110010000001"), ("0010110010000000"), ("0010110001111001"), ("0010110001110111"), ("0010110001110110"), ("0010110001110101"), ("0010110001110100"), ("0010110001110010"), ("0010110001110001"), ("0010110001110000"), ("0010110001101001"), ("0010110001100111"), ("0010110001100110"), ("0010110001100101"), ("0010110001100100"), ("0010110001100011"), ("0010110001100001"), ("0010110001100000"), ("0010110001011001"), ("0010110001011000"), ("0010110001010110"), ("0010110001010101"), ("0010110001010100"), ("0010110001010011"), ("0010110001010010"), ("0010110001010000"), ("0010110001001001"), ("0010110001001000"), ("0010110001000111"), ("0010110001000101"), ("0010110001000100"), ("0010110001000011"), ("0010110001000010"), ("0010110001000000"), ("0010110000111001"), ("0010110000111000"), ("0010110000110111"), ("0010110000110110"), ("0010110000110100"), ("0010110000110011"), ("0010110000110010"), ("0010110000110001"), ("0010110000101001"), ("0010110000101000"), ("0010110000100111"), ("0010110000100110"), ("0010110000100100"), ("0010110000100011"), ("0010110000100010"), ("0010110000100001"), ("0010110000011001"), ("0010110000011000"), ("0010110000010111"), ("0010110000010110"), ("0010110000010100"), ("0010110000010011"), ("0010110000010010"), ("0010110000010001"), ("0010110000001001"), ("0010110000001000"), ("0010110000000111"), ("0010110000000110"), ("0010110000000100"), ("0010110000000011"), ("0010110000000010"), ("0010110000000001"), ("0001110010011001"), ("0001110010011000"), ("0001110010010111"), ("0001110010010110"), ("0001110010010100"), ("0001110010010011"), ("0001110010010010"), ("0001110010010001"), ("0001110010001001"), ("0001110010001000"), ("0001110010000111"), ("0001110010000110"), ("0001110010000100"), ("0001110010000011"), ("0001110010000010"), ("0001110010000001"), ("0001110001111001"), ("0001110001111000"), ("0001110001110111"), ("0001110001110110"), ("0001110001110101"), ("0001110001110011"), ("0001110001110010"), ("0001110001110001"), ("0001110001110000"), ("0001110001101001"), ("0001110001100111"), ("0001110001100110"), ("0001110001100101"), ("0001110001100100"), ("0001110001100011"), ("0001110001100010"), ("0001110001100001"), ("0001110001100000"), ("0001110001011000"), ("0001110001010111"), ("0001110001010110"), ("0001110001010101"), ("0001110001010100"), ("0001110001010011"), ("0001110001010010"), ("0001110001010001"), ("0001110001010000"), ("0001110001001001"), ("0001110001001000"), ("0001110001000111"), ("0001110001000110"), ("0001110001000101"), ("0001110001000100"), ("0001110001000011"), ("0001110001000010"), ("0001110001000010"), ("0001110001000001"), ("0001110001000000"), ("0001110000111001"), ("0001110000111000"), ("0001110000111000"), ("0001110000110111"), ("0001110000110110"), ("0001110000110101"), ("0001110000110101"), ("0001110000110100"), ("0001110000110011"), ("0001110000110011"), ("0001110000110010"), ("0001110000110010"), ("0001110000110001"), ("0001110000110000"), ("0001110000110000"), ("0001110000101001"), ("0001110000101001"), ("0001110000101001"), ("0001110000101000"), ("0001110000101000"), ("0001110000101000"), ("0001110000100111"), ("0001110000100111"), ("0001110000100111"), ("0001110000100111"), ("0001110000100110"), ("0001110000100110"), ("0001110000100110"), ("0001110000100110"), ("0001110000100110"), ("0001110000100110"), ("0001110000100110"), ("0001110000100110"), ("0001110000100111"), ("0001110000100111"), ("0001110000100111"), ("0001110000100111"), ("0001110000100111"), ("0001110000101000"), ("0001110000101000"), ("0001110000101001"), ("0001110000101001"), ("0001110000110000"), ("0001110000110000"), ("0001110000110001"), ("0001110000110010"), ("0001110000110010"), ("0001110000110011"), ("0001110000110100"), ("0001110000110101"), ("0001110000110110"), ("0001110000110111"), ("0001110000111000"), ("0001110000111001"), ("0001110001000000"), ("0001110001000001"), ("0001110001000011"), ("0001110001000100"), ("0001110001000101"), ("0001110001000111"), ("0001110001001000"), ("0001110001010000"), ("0001110001010001"), ("0001110001010011"), ("0001110001010101"), ("0001110001010111"), ("0001110001011001"), ("0001110001100001"), ("0001110001100011"), ("0001110001100101"), ("0001110001100111"), ("0001110001101001"), ("0001110001110010"), ("0001110001110100"), ("0001110001110111"), ("0001110001111001"), ("0001110010000010"), ("0001110010000100"), ("0001110010000111"), ("0001110010010000"), ("0001110010010011"), ("0001110010010110"), ("0001110010011001"), ("0010110000000011"), ("0010110000000110"), ("0010110000001001"), ("0010110000010011"), ("0010110000010110"), ("0010110000100000"), ("0010110000100100"), ("0010110000101000"), ("0010110000110010"), ("0010110000110110"), ("0010110001000000"), ("0010110001000100"), ("0010110001001000"), ("0010110001010011"), ("0010110001010111"), ("0010110001100010"), ("0010110001100111"), ("0010110001110001"), ("0010110001110110"), ("0010110010000001"), ("0010110010000111"), ("0010110010010010"), ("0010110010010111"), ("0011110000000011"), ("0011110000001000"), ("0011110000010100"), ("0011110000100000"), ("0011110000100110"), ("0011110000110010"), ("0011110000111000"), ("0011110001000101"), ("0011110001010001"), ("0011110001011000"), ("0011110001100100"), ("0011110001110001"), ("0011110001111000"), ("0011110010000101"), ("0011110010010010"), ("0100110000000000"), ("0100110000000111"), ("0100110000010101"), ("0100110000100010"), ("0100110000110000"), ("0100110000111000"));

    begin
    -- Internal processes ----------------------------------------------------------
    select_rom : process(voltage, en_dists_cm, en_dists_in)
    begin
        if (en_dists_cm = '1') then
            distance <= dists_cm(CONV_INTEGER(UNSIGNED(voltage)));
        elsif (en_dists_in = '1') then
            distance <= dists_in(CONV_INTEGER(UNSIGNED(voltage)));
        else
            distance <= "1111" & "1111" & "1111" & "1111";
        end if;
    end process ; -- select_rom
    
end Behavioral;
    
