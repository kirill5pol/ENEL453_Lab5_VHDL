library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    use IEEE.STD_LOGIC_ARITH.ALL;
    use IEEE.STD_LOGIC_UNSIGNED.ALL;
    
    entity estimator is
            generic (width: integer := 9);
            Port (
                    clk        : in  STD_LOGIC;
                    reset      : in  STD_LOGIC;
                    en_dists_mm: in STD_LOGIC;
                    en_dists_cm: in STD_LOGIC;
                    en_dists_in: in STD_LOGIC;
                    voltage    : in  STD_LOGIC_VECTOR(width-1 downto 0);
                    distance   : out STD_LOGIC_VECTOR(3*4-1 downto 0)
            );
    end estimator;
    
    architecture Behavioral of estimator is
    type ROM is array (0 to 511) of STD_LOGIC_VECTOR(8 downto 0);
    constant dists_mm: ROM := (("011000100011"), ("011000010111"), ("011000010000"), ("011000000100"), ("010110010111"), ("010110010001"), ("010110000101"), ("010101111000"), ("010101110010"), ("010101100110"), ("010101100000"), ("010101010100"), ("010101001000"), ("010101000010"), ("010100110110"), ("010100110000"), ("010100100101"), ("010100011001"), ("010100010100"), ("010100001000"), ("010100000010"), ("010010010111"), ("010010010010"), ("010010000110"), ("010010000001"), ("010001110110"), ("010001110001"), ("010001100110"), ("010001100000"), ("010001010101"), ("010001010001"), ("010001000110"), ("010001000001"), ("010000110110"), ("010000110001"), ("010000100110"), ("010000100010"), ("010000010111"), ("010000010011"), ("010000001000"), ("010000000100"), ("001110011001"), ("001110010101"), ("001110010001"), ("001110000110"), ("001110000010"), ("001101111000"), ("001101110100"), ("001101110000"), ("001101100110"), ("001101100010"), ("001101011000"), ("001101010100"), ("001101010000"), ("001101000110"), ("001101000010"), ("001100111000"), ("001100110101"), ("001100110001"), ("001100101000"), ("001100100100"), ("001100100000"), ("001100010111"), ("001100010011"), ("001100010000"), ("001100000111"), ("001100000011"), ("001100000000"), ("001010010111"), ("001010010100"), ("001010010000"), ("001010000111"), ("001010000100"), ("001010000001"), ("001001111000"), ("001001110101"), ("001001110010"), ("001001101001"), ("001001100110"), ("001001100011"), ("001001100001"), ("001001011000"), ("001001010101"), ("001001010010"), ("001001010000"), ("001001000111"), ("001001000100"), ("001001000010"), ("001000111001"), ("001000110111"), ("001000110100"), ("001000110010"), ("001000101001"), ("001000100111"), ("001000100100"), ("001000100010"), ("001000100000"), ("001000011000"), ("001000010101"), ("001000010011"), ("001000010001"), ("001000001001"), ("001000000111"), ("001000000100"), ("001000000010"), ("001000000000"), ("000110011000"), ("000110010110"), ("000110010100"), ("000110010010"), ("000110010000"), ("000110001001"), ("000110000111"), ("000110000101"), ("000110000011"), ("000110000001"), ("000101111001"), ("000101111000"), ("000101110110"), ("000101110100"), ("000101110011"), ("000101110001"), ("000101101001"), ("000101101000"), ("000101100110"), ("000101100101"), ("000101100011"), ("000101100010"), ("000101100000"), ("000101011001"), ("000101010111"), ("000101010110"), ("000101010100"), ("000101010011"), ("000101010010"), ("000101010000"), ("000101001001"), ("000101001000"), ("000101000110"), ("000101000101"), ("000101000100"), ("000101000010"), ("000101000001"), ("000101000000"), ("000100111001"), ("000100111000"), ("000100110111"), ("000100110101"), ("000100110100"), ("000100110011"), ("000100110010"), ("000100110001"), ("000100110000"), ("000100101001"), ("000100101000"), ("000100100111"), ("000100100110"), ("000100100101"), ("000100100100"), ("000100100011"), ("000100100010"), ("000100100001"), ("000100100000"), ("000100100000"), ("000100011001"), ("000100011000"), ("000100010111"), ("000100010110"), ("000100010101"), ("000100010100"), ("000100010100"), ("000100010011"), ("000100010010"), ("000100010001"), ("000100010001"), ("000100010000"), ("000100001001"), ("000100001000"), ("000100001000"), ("000100000111"), ("000100000110"), ("000100000110"), ("000100000101"), ("000100000100"), ("000100000100"), ("000100000011"), ("000100000011"), ("000100000010"), ("000100000001"), ("000100000001"), ("000100000000"), ("000100000000"), ("100110010101"), ("100110010000"), ("100110000100"), ("100101111001"), ("100101110100"), ("100101101000"), ("100101100011"), ("100101011000"), ("100101010011"), ("100101001000"), ("100101000011"), ("100100111001"), ("100100110100"), ("100100101001"), ("100100100101"), ("100100100000"), ("100100010110"), ("100100010010"), ("100100000111"), ("100100000011"), ("100010011001"), ("100010010101"), ("100010010001"), ("100010000111"), ("100010000011"), ("100001111001"), ("100001110101"), ("100001110001"), ("100001101000"), ("100001100100"), ("100001100000"), ("100001010111"), ("100001010011"), ("100001010000"), ("100001000110"), ("100001000011"), ("100001000000"), ("100000110110"), ("100000110011"), ("100000110000"), ("100000100110"), ("100000100011"), ("100000100000"), ("100000010111"), ("100000010100"), ("100000010001"), ("100000001000"), ("100000000101"), ("100000000010"), ("011110011001"), ("011110010110"), ("011110010011"), ("011110010000"), ("011110000111"), ("011110000100"), ("011110000010"), ("011101111001"), ("011101110110"), ("011101110011"), ("011101110001"), ("011101101000"), ("011101100101"), ("011101100011"), ("011101100000"), ("011101010111"), ("011101010101"), ("011101010010"), ("011101010000"), ("011101000111"), ("011101000100"), ("011101000010"), ("011100111001"), ("011100110111"), ("011100110100"), ("011100110010"), ("011100101001"), ("011100100111"), ("011100100100"), ("011100100010"), ("011100011001"), ("011100010111"), ("011100010100"), ("011100010010"), ("011100001001"), ("011100000111"), ("011100000101"), ("011100000010"), ("011100000000"), ("011010010111"), ("011010010101"), ("011010010010"), ("011010010000"), ("011010001000"), ("011010000101"), ("011010000011"), ("011010000000"), ("011001111000"), ("011001110101"), ("011001110011"), ("011001110001"), ("011001101000"), ("011001100110"), ("011001100011"), ("011001100001"), ("011001011000"), ("011001010110"), ("011001010100"), ("011001010001"), ("011001001001"), ("011001000110"), ("011001000100"), ("011001000001"), ("011000111001"), ("011000110110"), ("011000110100"), ("011000110001"), ("011000101001"), ("011000100111"), ("011000100100"), ("011000100010"), ("011000011001"), ("011000010111"), ("011000010100"), ("011000010010"), ("011000001001"), ("011000000111"), ("011000000100"), ("011000000010"), ("010110011001"), ("010110010111"), ("010110010100"), ("010110010010"), ("010110001001"), ("010110000111"), ("010110000100"), ("010110000010"), ("010101111001"), ("010101110111"), ("010101110100"), ("010101110010"), ("010101101001"), ("010101100111"), ("010101100100"), ("010101100010"), ("010101011001"), ("010101010111"), ("010101010101"), ("010101010010"), ("010101010000"), ("010101000111"), ("010101000101"), ("010101000010"), ("010101000000"), ("010100110111"), ("010100110101"), ("010100110010"), ("010100110000"), ("010100101000"), ("010100100101"), ("010100100011"), ("010100100000"), ("010100011000"), ("010100010110"), ("010100010011"), ("010100010001"), ("010100001001"), ("010100000110"), ("010100000100"), ("010100000010"), ("010100000000"), ("010010010111"), ("010010010101"), ("010010010011"), ("010010010001"), ("010010001001"), ("010010000111"), ("010010000100"), ("010010000010"), ("010010000000"), ("010001111000"), ("010001110110"), ("010001110100"), ("010001110010"), ("010001110000"), ("010001101000"), ("010001100110"), ("010001100101"), ("010001100011"), ("010001100001"), ("010001011001"), ("010001010111"), ("010001010110"), ("010001010100"), ("010001010011"), ("010001010001"), ("010001001001"), ("010001001000"), ("010001000110"), ("010001000101"), ("010001000100"), ("010001000010"), ("010001000001"), ("010001000000"), ("010000111001"), ("010000110111"), ("010000110110"), ("010000110101"), ("010000110100"), ("010000110011"), ("010000110011"), ("010000110010"), ("010000110001"), ("010000110000"), ("010000110000"), ("010000101001"), ("010000101001"), ("010000101000"), ("010000101000"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000101000"), ("010000101000"), ("010000101000"), ("010000101001"), ("010000110000"), ("010000110000"), ("010000110001"), ("010000110010"), ("010000110011"), ("010000110100"), ("010000110101"), ("010000110110"), ("010000111000"), ("010000111001"), ("010001000001"), ("010001000010"), ("010001000100"), ("010001000110"), ("010001001000"), ("010001010000"), ("010001010010"), ("010001010100"), ("010001010111"), ("010001011001"), ("010001100010"), ("010001100101"), ("010001101000"), ("010001110001"), ("010001110100"), ("010001110111"), ("010010000000"), ("010010000100"), ("010010001000"), ("010010010001"), ("010010010101"), ("010010011001"), ("010100000100"), ("010100001000"), ("010100010010"), ("010100010111"), ("010100100010"), ("010100100111"), ("010100110010"), ("010100110111"), ("010101000010"), ("010101001000"), ("010101010100"), ("010101100000"), ("010101100110"), ("010101110010"), ("010101111000"), ("010110000101"), ("010110010010"), ("010110011000"), ("011000000110"), ("011000010011"), ("011000100000"), ("011000101000"), ("011000110110"), ("011001000100"), ("011001010010"), ("011001100000"), ("011001101001"), ("011001111000"), ("011010000111"), ("011010010110"), ("011100000101"), ("011100010101"), ("011100100101"), ("011100110101"), ("011101000101"), ("011101010110"), ("011101100110"), ("011101110111"), ("011110001000"), ("100000000000"), ("100000010001"), ("100000100011"), ("100000110101"), ("100001000111"), ("100001100000"), ("100001110011"), ("100010000110"), ("100010011001"), ("100100010010"), ("100100100110"), ("100101000000"), ("100101010101"), ("100101101001"), ("100110000100"), ("100110011001"), ("000100000001"), ("000100000011"), ("000100000100"));
    constant dists_cm: ROM := (("011000100011"), ("011000010111"), ("011000010000"), ("011000000100"), ("010110010111"), ("010110010001"), ("010110000101"), ("010101111000"), ("010101110010"), ("010101100110"), ("010101100000"), ("010101010100"), ("010101001000"), ("010101000010"), ("010100110110"), ("010100110000"), ("010100100101"), ("010100011001"), ("010100010100"), ("010100001000"), ("010100000010"), ("010010010111"), ("010010010010"), ("010010000110"), ("010010000001"), ("010001110110"), ("010001110001"), ("010001100110"), ("010001100000"), ("010001010101"), ("010001010001"), ("010001000110"), ("010001000001"), ("010000110110"), ("010000110001"), ("010000100110"), ("010000100010"), ("010000010111"), ("010000010011"), ("010000001000"), ("010000000100"), ("001110011001"), ("001110010101"), ("001110010001"), ("001110000110"), ("001110000010"), ("001101111000"), ("001101110100"), ("001101110000"), ("001101100110"), ("001101100010"), ("001101011000"), ("001101010100"), ("001101010000"), ("001101000110"), ("001101000010"), ("001100111000"), ("001100110101"), ("001100110001"), ("001100101000"), ("001100100100"), ("001100100000"), ("001100010111"), ("001100010011"), ("001100010000"), ("001100000111"), ("001100000011"), ("001100000000"), ("001010010111"), ("001010010100"), ("001010010000"), ("001010000111"), ("001010000100"), ("001010000001"), ("001001111000"), ("001001110101"), ("001001110010"), ("001001101001"), ("001001100110"), ("001001100011"), ("001001100001"), ("001001011000"), ("001001010101"), ("001001010010"), ("001001010000"), ("001001000111"), ("001001000100"), ("001001000010"), ("001000111001"), ("001000110111"), ("001000110100"), ("001000110010"), ("001000101001"), ("001000100111"), ("001000100100"), ("001000100010"), ("001000100000"), ("001000011000"), ("001000010101"), ("001000010011"), ("001000010001"), ("001000001001"), ("001000000111"), ("001000000100"), ("001000000010"), ("001000000000"), ("000110011000"), ("000110010110"), ("000110010100"), ("000110010010"), ("000110010000"), ("000110001001"), ("000110000111"), ("000110000101"), ("000110000011"), ("000110000001"), ("000101111001"), ("000101111000"), ("000101110110"), ("000101110100"), ("000101110011"), ("000101110001"), ("000101101001"), ("000101101000"), ("000101100110"), ("000101100101"), ("000101100011"), ("000101100010"), ("000101100000"), ("000101011001"), ("000101010111"), ("000101010110"), ("000101010100"), ("000101010011"), ("000101010010"), ("000101010000"), ("000101001001"), ("000101001000"), ("000101000110"), ("000101000101"), ("000101000100"), ("000101000010"), ("000101000001"), ("000101000000"), ("000100111001"), ("000100111000"), ("000100110111"), ("000100110101"), ("000100110100"), ("000100110011"), ("000100110010"), ("000100110001"), ("000100110000"), ("000100101001"), ("000100101000"), ("000100100111"), ("000100100110"), ("000100100101"), ("000100100100"), ("000100100011"), ("000100100010"), ("000100100001"), ("000100100000"), ("000100100000"), ("000100011001"), ("000100011000"), ("000100010111"), ("000100010110"), ("000100010101"), ("000100010100"), ("000100010100"), ("000100010011"), ("000100010010"), ("000100010001"), ("000100010001"), ("000100010000"), ("000100001001"), ("000100001000"), ("000100001000"), ("000100000111"), ("000100000110"), ("000100000110"), ("000100000101"), ("000100000100"), ("000100000100"), ("000100000011"), ("000100000011"), ("000100000010"), ("000100000001"), ("000100000001"), ("000100000000"), ("000100000000"), ("100110010101"), ("100110010000"), ("100110000100"), ("100101111001"), ("100101110100"), ("100101101000"), ("100101100011"), ("100101011000"), ("100101010011"), ("100101001000"), ("100101000011"), ("100100111001"), ("100100110100"), ("100100101001"), ("100100100101"), ("100100100000"), ("100100010110"), ("100100010010"), ("100100000111"), ("100100000011"), ("100010011001"), ("100010010101"), ("100010010001"), ("100010000111"), ("100010000011"), ("100001111001"), ("100001110101"), ("100001110001"), ("100001101000"), ("100001100100"), ("100001100000"), ("100001010111"), ("100001010011"), ("100001010000"), ("100001000110"), ("100001000011"), ("100001000000"), ("100000110110"), ("100000110011"), ("100000110000"), ("100000100110"), ("100000100011"), ("100000100000"), ("100000010111"), ("100000010100"), ("100000010001"), ("100000001000"), ("100000000101"), ("100000000010"), ("011110011001"), ("011110010110"), ("011110010011"), ("011110010000"), ("011110000111"), ("011110000100"), ("011110000010"), ("011101111001"), ("011101110110"), ("011101110011"), ("011101110001"), ("011101101000"), ("011101100101"), ("011101100011"), ("011101100000"), ("011101010111"), ("011101010101"), ("011101010010"), ("011101010000"), ("011101000111"), ("011101000100"), ("011101000010"), ("011100111001"), ("011100110111"), ("011100110100"), ("011100110010"), ("011100101001"), ("011100100111"), ("011100100100"), ("011100100010"), ("011100011001"), ("011100010111"), ("011100010100"), ("011100010010"), ("011100001001"), ("011100000111"), ("011100000101"), ("011100000010"), ("011100000000"), ("011010010111"), ("011010010101"), ("011010010010"), ("011010010000"), ("011010001000"), ("011010000101"), ("011010000011"), ("011010000000"), ("011001111000"), ("011001110101"), ("011001110011"), ("011001110001"), ("011001101000"), ("011001100110"), ("011001100011"), ("011001100001"), ("011001011000"), ("011001010110"), ("011001010100"), ("011001010001"), ("011001001001"), ("011001000110"), ("011001000100"), ("011001000001"), ("011000111001"), ("011000110110"), ("011000110100"), ("011000110001"), ("011000101001"), ("011000100111"), ("011000100100"), ("011000100010"), ("011000011001"), ("011000010111"), ("011000010100"), ("011000010010"), ("011000001001"), ("011000000111"), ("011000000100"), ("011000000010"), ("010110011001"), ("010110010111"), ("010110010100"), ("010110010010"), ("010110001001"), ("010110000111"), ("010110000100"), ("010110000010"), ("010101111001"), ("010101110111"), ("010101110100"), ("010101110010"), ("010101101001"), ("010101100111"), ("010101100100"), ("010101100010"), ("010101011001"), ("010101010111"), ("010101010101"), ("010101010010"), ("010101010000"), ("010101000111"), ("010101000101"), ("010101000010"), ("010101000000"), ("010100110111"), ("010100110101"), ("010100110010"), ("010100110000"), ("010100101000"), ("010100100101"), ("010100100011"), ("010100100000"), ("010100011000"), ("010100010110"), ("010100010011"), ("010100010001"), ("010100001001"), ("010100000110"), ("010100000100"), ("010100000010"), ("010100000000"), ("010010010111"), ("010010010101"), ("010010010011"), ("010010010001"), ("010010001001"), ("010010000111"), ("010010000100"), ("010010000010"), ("010010000000"), ("010001111000"), ("010001110110"), ("010001110100"), ("010001110010"), ("010001110000"), ("010001101000"), ("010001100110"), ("010001100101"), ("010001100011"), ("010001100001"), ("010001011001"), ("010001010111"), ("010001010110"), ("010001010100"), ("010001010011"), ("010001010001"), ("010001001001"), ("010001001000"), ("010001000110"), ("010001000101"), ("010001000100"), ("010001000010"), ("010001000001"), ("010001000000"), ("010000111001"), ("010000110111"), ("010000110110"), ("010000110101"), ("010000110100"), ("010000110011"), ("010000110011"), ("010000110010"), ("010000110001"), ("010000110000"), ("010000110000"), ("010000101001"), ("010000101001"), ("010000101000"), ("010000101000"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000100111"), ("010000101000"), ("010000101000"), ("010000101000"), ("010000101001"), ("010000110000"), ("010000110000"), ("010000110001"), ("010000110010"), ("010000110011"), ("010000110100"), ("010000110101"), ("010000110110"), ("010000111000"), ("010000111001"), ("010001000001"), ("010001000010"), ("010001000100"), ("010001000110"), ("010001001000"), ("010001010000"), ("010001010010"), ("010001010100"), ("010001010111"), ("010001011001"), ("010001100010"), ("010001100101"), ("010001101000"), ("010001110001"), ("010001110100"), ("010001110111"), ("010010000000"), ("010010000100"), ("010010001000"), ("010010010001"), ("010010010101"), ("010010011001"), ("010100000100"), ("010100001000"), ("010100010010"), ("010100010111"), ("010100100010"), ("010100100111"), ("010100110010"), ("010100110111"), ("010101000010"), ("010101001000"), ("010101010100"), ("010101100000"), ("010101100110"), ("010101110010"), ("010101111000"), ("010110000101"), ("010110010010"), ("010110011000"), ("011000000110"), ("011000010011"), ("011000100000"), ("011000101000"), ("011000110110"), ("011001000100"), ("011001010010"), ("011001100000"), ("011001101001"), ("011001111000"), ("011010000111"), ("011010010110"), ("011100000101"), ("011100010101"), ("011100100101"), ("011100110101"), ("011101000101"), ("011101010110"), ("011101100110"), ("011101110111"), ("011110001000"), ("100000000000"), ("100000010001"), ("100000100011"), ("100000110101"), ("100001000111"), ("100001100000"), ("100001110011"), ("100010000110"), ("100010011001"), ("100100010010"), ("100100100110"), ("100101000000"), ("100101010101"), ("100101101001"), ("100110000100"), ("100110011001"), ("000100000001"), ("000100000011"), ("000100000100"));
    constant dists_in: ROM := (("001001000101"), ("001001000010"), ("001001000000"), ("001000110111"), ("001000110101"), ("001000110010"), ("001000110000"), ("001000100111"), ("001000100101"), ("001000100011"), ("001000100000"), ("001000011000"), ("001000010101"), ("001000010011"), ("001000010001"), ("001000001001"), ("001000000110"), ("001000000100"), ("001000000010"), ("001000000000"), ("000110011000"), ("000110010101"), ("000110010011"), ("000110010001"), ("000110001001"), ("000110000111"), ("000110000101"), ("000110000011"), ("000110000001"), ("000101111001"), ("000101110111"), ("000101110101"), ("000101110011"), ("000101110001"), ("000101101001"), ("000101101000"), ("000101100110"), ("000101100100"), ("000101100010"), ("000101100000"), ("000101011001"), ("000101010111"), ("000101010101"), ("000101010011"), ("000101010010"), ("000101010000"), ("000101001000"), ("000101000111"), ("000101000101"), ("000101000100"), ("000101000010"), ("000101000000"), ("000100111001"), ("000100110111"), ("000100110110"), ("000100110100"), ("000100110011"), ("000100110010"), ("000100110000"), ("000100101001"), ("000100100111"), ("000100100110"), ("000100100100"), ("000100100011"), ("000100100010"), ("000100100000"), ("000100011001"), ("000100011000"), ("000100010111"), ("000100010101"), ("000100010100"), ("000100010011"), ("000100010010"), ("000100010000"), ("000100001001"), ("000100001000"), ("000100000111"), ("000100000110"), ("000100000100"), ("000100000011"), ("000100000010"), ("000100000001"), ("000100000000"), ("100110010101"), ("100110000100"), ("100101110100"), ("100101100011"), ("100101010011"), ("100101000011"), ("100100110011"), ("100100100011"), ("100100010011"), ("100100000100"), ("100010010100"), ("100010000101"), ("100001110110"), ("100001100111"), ("100001011000"), ("100001001001"), ("100001000000"), ("100000110010"), ("100000100011"), ("100000010101"), ("100000000110"), ("011110011000"), ("011110010000"), ("011110000010"), ("011101110100"), ("011101100110"), ("011101011001"), ("011101010001"), ("011101000100"), ("011100110110"), ("011100101001"), ("011100100010"), ("011100010101"), ("011100001000"), ("011100000001"), ("011010010100"), ("011010001000"), ("011010000001"), ("011001110101"), ("011001101000"), ("011001100010"), ("011001010110"), ("011001001001"), ("011001000011"), ("011000110111"), ("011000110010"), ("011000100110"), ("011000100000"), ("011000010100"), ("011000001001"), ("011000000011"), ("010110011000"), ("010110010011"), ("010110000111"), ("010110000010"), ("010101110111"), ("010101110010"), ("010101100111"), ("010101100010"), ("010101011000"), ("010101010011"), ("010101001000"), ("010101000100"), ("010100111001"), ("010100110101"), ("010100110000"), ("010100100110"), ("010100100010"), ("010100010111"), ("010100010011"), ("010100001001"), ("010100000101"), ("010100000001"), ("010010010111"), ("010010010100"), ("010010010000"), ("010010000110"), ("010010000011"), ("010001111001"), ("010001110101"), ("010001110010"), ("010001101001"), ("010001100101"), ("010001100010"), ("010001011001"), ("010001010101"), ("010001010010"), ("010001001001"), ("010001000110"), ("010001000011"), ("010001000000"), ("010000110111"), ("010000110100"), ("010000110001"), ("010000101001"), ("010000100110"), ("010000100011"), ("010000100000"), ("010000011000"), ("010000010101"), ("010000010011"), ("010000010000"), ("010000001000"), ("010000000101"), ("010000000011"), ("010000000001"), ("001110011000"), ("001110010110"), ("001110010100"), ("001110010001"), ("001110001001"), ("001110000111"), ("001110000101"), ("001110000011"), ("001110000001"), ("001101111001"), ("001101110111"), ("001101110101"), ("001101110011"), ("001101110001"), ("001101101001"), ("001101100111"), ("001101100110"), ("001101100100"), ("001101100010"), ("001101100000"), ("001101011001"), ("001101010111"), ("001101010101"), ("001101010100"), ("001101010010"), ("001101010000"), ("001101001001"), ("001101000111"), ("001101000110"), ("001101000100"), ("001101000011"), ("001101000001"), ("001101000000"), ("001100111000"), ("001100110111"), ("001100110110"), ("001100110100"), ("001100110011"), ("001100110010"), ("001100110000"), ("001100101001"), ("001100101000"), ("001100100110"), ("001100100101"), ("001100100100"), ("001100100011"), ("001100100001"), ("001100100000"), ("001100011001"), ("001100011000"), ("001100010111"), ("001100010101"), ("001100010100"), ("001100010011"), ("001100010010"), ("001100010001"), ("001100010000"), ("001100001001"), ("001100000111"), ("001100000110"), ("001100000101"), ("001100000100"), ("001100000011"), ("001100000010"), ("001100000001"), ("001100000000"), ("001010011001"), ("001010011000"), ("001010010111"), ("001010010110"), ("001010010101"), ("001010010100"), ("001010010011"), ("001010010010"), ("001010010001"), ("001010010000"), ("001010001001"), ("001010001000"), ("001010000111"), ("001010000110"), ("001010000101"), ("001010000100"), ("001010000011"), ("001010000010"), ("001010000001"), ("001010000000"), ("001001111001"), ("001001111000"), ("001001110111"), ("001001110110"), ("001001110101"), ("001001110100"), ("001001110011"), ("001001110010"), ("001001110001"), ("001001110000"), ("001001101001"), ("001001101000"), ("001001101000"), ("001001100111"), ("001001100110"), ("001001100101"), ("001001100100"), ("001001100011"), ("001001100010"), ("001001100001"), ("001001100000"), ("001001011001"), ("001001011000"), ("001001010111"), ("001001010110"), ("001001010101"), ("001001010100"), ("001001010011"), ("001001010010"), ("001001010001"), ("001001010000"), ("001001001001"), ("001001001000"), ("001001000111"), ("001001000110"), ("001001000101"), ("001001000100"), ("001001000011"), ("001001000010"), ("001001000010"), ("001001000001"), ("001001000000"), ("001000111001"), ("001000111000"), ("001000110111"), ("001000110110"), ("001000110101"), ("001000110100"), ("001000110011"), ("001000110010"), ("001000110001"), ("001000110000"), ("001000101001"), ("001000101000"), ("001000100111"), ("001000100110"), ("001000100101"), ("001000100100"), ("001000100011"), ("001000100010"), ("001000100001"), ("001000100000"), ("001000011001"), ("001000011000"), ("001000010111"), ("001000010110"), ("001000010101"), ("001000010100"), ("001000010011"), ("001000010010"), ("001000010001"), ("001000010000"), ("001000001001"), ("001000001000"), ("001000000111"), ("001000000110"), ("001000000110"), ("001000000101"), ("001000000100"), ("001000000011"), ("001000000010"), ("001000000001"), ("001000000000"), ("000110011001"), ("000110011000"), ("000110010111"), ("000110010110"), ("000110010110"), ("000110010101"), ("000110010100"), ("000110010011"), ("000110010010"), ("000110010001"), ("000110010000"), ("000110010000"), ("000110001001"), ("000110001000"), ("000110000111"), ("000110000110"), ("000110000110"), ("000110000101"), ("000110000100"), ("000110000011"), ("000110000011"), ("000110000010"), ("000110000001"), ("000110000000"), ("000110000000"), ("000101111001"), ("000101111000"), ("000101111000"), ("000101110111"), ("000101110111"), ("000101110110"), ("000101110101"), ("000101110101"), ("000101110100"), ("000101110100"), ("000101110011"), ("000101110011"), ("000101110010"), ("000101110010"), ("000101110010"), ("000101110001"), ("000101110001"), ("000101110000"), ("000101110000"), ("000101110000"), ("000101101001"), ("000101101001"), ("000101101001"), ("000101101001"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101000"), ("000101101001"), ("000101101001"), ("000101101001"), ("000101101001"), ("000101110000"), ("000101110000"), ("000101110001"), ("000101110001"), ("000101110001"), ("000101110010"), ("000101110011"), ("000101110011"), ("000101110100"), ("000101110100"), ("000101110101"), ("000101110110"), ("000101110111"), ("000101111000"), ("000101111001"), ("000110000000"), ("000110000001"), ("000110000010"), ("000110000011"), ("000110000100"), ("000110000101"), ("000110000110"), ("000110000111"), ("000110001001"), ("000110010000"), ("000110010010"), ("000110010011"), ("000110010101"), ("000110010110"), ("000110011000"), ("001000000000"), ("001000000001"), ("001000000011"), ("001000000101"), ("001000000111"), ("001000001001"), ("001000010001"), ("001000010011"), ("001000010101"), ("001000011000"), ("001000100000"), ("001000100010"), ("001000100101"), ("001000100111"), ("001000110000"), ("001000110011"), ("001000110101"), ("001000111000"), ("001001000001"), ("001001000100"), ("001001000111"), ("001001010000"), ("001001010011"), ("001001010110"), ("001001100000"), ("001001100011"), ("001001100111"), ("001001110000"), ("001001110100"), ("001001110111"), ("001010000001"), ("001010000101"), ("001010001001"), ("001010010011"), ("001010010111"), ("001100000001"), ("001100000110"), ("001100010000"), ("001100010100"), ("001100011001"), ("001100100100"), ("001100101000"), ("001100110011"), ("001100111000"), ("001101000011"), ("001101001000"), ("001101010100"), ("001101011001"), ("001101100100"), ("001101110000"), ("001101110110"), ("001110000001"), ("001110000111"), ("001110010011"), ("001110011001"), ("010000000101"), ("010000010001"));

    begin
    -- Internal processes ----------------------------------------------------------
    select_rom : process(en_dists_mm,  en_dists_cm,  en_dists_in)
    begin
        if (en_dists_mm = '1') then
            distance <= dists_mm(CONV_INTEGER(UNSIGNED(voltage)));
        elsif (en_dists_cm = '1') then
            distance <= dists_cm(CONV_INTEGER(UNSIGNED(voltage)));
        elsif (en_dists_in = '1') then
            distance <= dists_in(CONV_INTEGER(UNSIGNED(voltage)));
        else
            distance <= "1111" & "1111" & "1111";
        end if;
    end process ; -- select_rom
    
end Behavioral;
    
