--
--    Digits Box: takes in 3 digits (from 0 to 9) and prints those digits on the 
--                vga monitor.
--    
--    Module of:
--        - vga_module
--
--    Internal singals:
--        - sig_0 - sig_10: A 5x5 matrix that contains a digit from 0-9
--        - sig_dec: A matrix the contains an image of a decimal point
--        - box_loc_x/y_min/max: Min and max indices from x and y
--        - pixel_color: Colour of an individual pixel


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity digits_box is
    Port ( 	clk : in  STD_LOGIC;
			reset : in  STD_LOGIC;

            digit_tens: in STD_LOGIC_VECTOR(3 downto 0); -- Max number is 9 so we need 4 bits
            digit_ones: in STD_LOGIC_VECTOR(3 downto 0); -- Max number is 9 so we need 4 bits
            digit_tenths: in STD_LOGIC_VECTOR(3 downto 0); -- Max number is 9 so we need 4 bits

			scan_line_x: in STD_LOGIC_VECTOR(10 downto 0);
			scan_line_y: in STD_LOGIC_VECTOR(10 downto 0);
			kHz: in STD_LOGIC;
			red: out STD_LOGIC_VECTOR(3 downto 0);
			blue: out STD_LOGIC_VECTOR(3 downto 0);
			green: out std_logic_vector(3 downto 0)
		  );
end digits_box;

architecture Behavioral of digits_box is

-- Internal Signals  -----------------------------------------------------------
    -- You have 3 digits + 1 decimal point -> 50 by 50 for each -> width 200, height 50
    type MAT is array (24 downto 0) of std_logic_vector(24 downto 0);
    constant sig_0: MAT := (("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"));
    constant sig_1: MAT := (("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"));
    constant sig_2: MAT := (("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"));
    constant sig_3: MAT := (("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"));
    constant sig_4: MAT := (("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("0000011111000001111100000"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"));
    constant sig_5: MAT := (("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000111111111100000"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("0000000000000000000011111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"));
    constant sig_6: MAT := (("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111111111111111111100000"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"));
    constant sig_7: MAT := (("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("1111111111111111111111111"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000000000111110000000000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("0000011111000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"), ("1111100000000000000000000"));
    constant sig_8: MAT := (("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"), ("0000011111111111111100000"));
    constant sig_9: MAT := (("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("1111100000000000000011111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000011111111111111111111"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("0000000000000001111100000"), ("1111111111111110000000000"), ("1111111111111110000000000"), ("1111111111111110000000000"), ("1111111111111110000000000"), ("1111111111111110000000000"));

    constant box_loc_x_min: std_logic_vector(9 downto 0) := "0000000000";
    constant box_loc_y_min: std_logic_vector(9 downto 0) := "0000000000";
    constant box_loc_x_max: std_logic_vector(9 downto 0) := "1001111111"; -- 640-1 -- 640 is 1010000000
    constant box_loc_y_max: std_logic_vector(9 downto 0) := "0111011111"; -- 480-1 -- 480 is 0111100000
    signal pixel_color: std_logic_vector(11 downto 0);

    -- Offset from 0,0 for digits & scale factor
    constant offset_x: STD_LOGIC_VECTOR(9 downto 0) := "0000010000"; -- Offset 16 pixels
    constant offset_y: STD_LOGIC_VECTOR(9 downto 0) := "0000010000"; -- Offset 16 pixels
    constant digit_size: STD_LOGIC_VECTOR(6 downto 0) := "0011001"; -- Max size of a digit is 127x127
begin

-- Internal processes  ---------------------------------------------------------
    pixel_color <= "111111111111"; -- TODO make this work...
    --pixel_color <= ( -- When it matches a pixel representing a digit
    --                    (  
    --                        box_color AND 
    --                        initials(index_of_initials)
    --                    ) OR 
    --                    (
    --                        "111111111111" AND 
    --                        (NOT initials(index_of_initials)))
    --                    ) 
    --          when  ((scan_line_x >= box_loc_x) and 
    --                 (scan_line_y >= box_loc_y) and 
    --                 (scan_line_x < box_loc_x+box_width) and 
    --                 (scan_line_y < box_loc_y+box_width))
    --        else
    --                 "111111111111"; -- represents WHITE
								
red   <= pixel_color(11 downto 8);
green <= pixel_color(7 downto 4);
blue  <= pixel_color(3 downto 0);


end Behavioral;

